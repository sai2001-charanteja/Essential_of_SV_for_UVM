class sequencer extends component_base;
	
	
	function new(string name,component_base parent);
		super.new(name,parent);
	endfunction
	
endclass
