package packet_pkg;
	
	`include "packet_data.sv"

endpackage